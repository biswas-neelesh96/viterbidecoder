
module viterbi_decoder(input [1:0]dec_in,
                       input [1:0]w0_000,w0_001,w1_010,w1_011,w2_100,w2_101,w3_110,w3_111,
                       input [1:0]w4_000,w4_001,w5_010,w5_011,w6_100,w6_101,w7_110,w7_111,
                       input clk,sel0,rst,
                       input [1:0]sel1, 
                       
                       output [2:0]s0_000,s0_001,s1_010,s1_011,s2_100,s2_101,s3_110,s3_111,
                       output [2:0]s4_000,s4_001,s5_010,s5_011,s6_100,s6_101,s7_110,s7_111,
                       output [2:0]r000,r001,r010,r011,r100,r101,r110,r111,
                       output [2:0]out);
//wire [1:0]s0_00,s0_01,s1_10,s1_11,s2_00,s2_01,s3_10,s3_11;
//wire [1:0]r00,r01,r10,r11;
    
bmu b0 (dec_in,w0_000,w0_001,w1_010,w1_011,w2_100,w2_101,w3_110,w3_111,w4_000,w4_001,w5_010,w5_011,w6_100,w6_101,w7_110,w7_111,
               s0_000,s0_001,s1_010,s1_011,s2_100,s2_101,s3_110,s3_111,s4_000,s4_001,s5_010,s5_011,s6_100,s6_101,s7_110,s7_111);
pmu p0 ( s0_000,s0_001,s1_010,s1_011,s2_100,s2_101,s3_110,s3_111,s4_000,s4_001,s5_010,s5_011,s6_100,s6_101,s7_110,s7_111,clk,sel0,rst,sel1,r000,r001,r010,r011,r100,r101,r110,r111);
smu s0 (r000,r001,r010,r011,r100,r101,r110,r111,clk,rst,out);

endmodule